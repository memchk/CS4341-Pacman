module dummy;
endmodule