module map_ram (
    input logic i_clk, i_write, i_en,
    input logic [5:0] i_tile_x,
    input logic [4:0] i_tile_y,
    output logic o_tile_value
);

reg [49:0] r_map_ram [32];

initial begin
    r_map_ram[00] = 50'b11111111111111111111111111111111111111111111111111;
    r_map_ram[01] = 50'b10000000000001111000000000010000000000000000000001;
    r_map_ram[02] = 50'b10111111111101111011111111011111111110000000000101;
    r_map_ram[03] = 50'b10100000000101100010000001010000000010000000000101;
    r_map_ram[04] = 50'b10111111111101101110000001010000000010000000000101;
    r_map_ram[05] = 50'b10000000000001101000000001010000000010000000000101;
    r_map_ram[06] = 50'b10111111111101101111111111011111111110111111111101;
    r_map_ram[07] = 50'b10100000000101100000000000000000000000000000000001;
    r_map_ram[08] = 50'b10111111111101101111111111111111111111111111111101;
    r_map_ram[09] = 50'b00000000000000001000000000000000000000000000000100;
    r_map_ram[10] = 50'b10000011000000001000000000000000000000000000000101;
    r_map_ram[11] = 50'b10000011000000000000000000000000000000000000000101;
    r_map_ram[12] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[13] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[14] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[15] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[16] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[17] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[18] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[19] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[20] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[21] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[22] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[23] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[24] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[25] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[26] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[27] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[28] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[29] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[30] = 50'b10000011000000000000000000000000000000000000000001;
    r_map_ram[31] = 50'b11111111111111111111111111111111111111111111111111;
end

always_ff @(posedge i_clk) begin
    if(i_en) begin
        if(i_write) begin
            r_map_ram[i_tile_y][i_tile_x] <= '0;
        end else begin
            o_tile_value <= r_map_ram[i_tile_y][i_tile_x];
        end
    end
end

endmodule