`default_nettype none